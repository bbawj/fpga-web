module mdio(
  input clk;
  );

  always @(posedge clk) begin
  end

endmodule
